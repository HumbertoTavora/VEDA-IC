module GPINAND(I0,I1,I2,I3,paridade_par);

input wire I0;
input wire I1;
input wire I2;
input wire I3;
output wire paridade_par;

wire	SYNTHESIZED_WIRE_09;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;

assign	SYNTHESIZED_WIRE_09 = ~(I0 & I0);

assign	SYNTHESIZED_WIRE_10 = ~(I1 & I1);

assign	SYNTHESIZED_WIRE_11 = ~(I2 & I2);

assign	SYNTHESIZED_WIRE_12 = ~(I3 & I3);

assign	SYNTHESIZED_WIRE_13 = ~(SYNTHESIZED_WIRE_09 & I1);

assign	SYNTHESIZED_WIRE_14 = ~(I0 & SYNTHESIZED_WIRE_10);

assign	SYNTHESIZED_WIRE_15 = ~(SYNTHESIZED_WIRE_11 & I3);

assign	SYNTHESIZED_WIRE_16 = ~(I2 & SYNTHESIZED_WIRE_12);

assign	SYNTHESIZED_WIRE_17 = ~(SYNTHESIZED_WIRE_13 & SYNTHESIZED_WIRE_14);

assign	SYNTHESIZED_WIRE_18 = ~(SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_16);

assign	SYNTHESIZED_WIRE_21 = ~(SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_17);

assign	SYNTHESIZED_WIRE_22 = ~(SYNTHESIZED_WIRE_18 & SYNTHESIZED_WIRE_18);

assign	SYNTHESIZED_WIRE_25 = ~(SYNTHESIZED_WIRE_21 & SYNTHESIZED_WIRE_18);

assign	SYNTHESIZED_WIRE_26 = ~(SYNTHESIZED_WIRE_22 & SYNTHESIZED_WIRE_17);

assign	paridade_par = ~(SYNTHESIZED_WIRE_25 & SYNTHESIZED_WIRE_26);


endmodule